module keyboard_testbech();

endmodule
